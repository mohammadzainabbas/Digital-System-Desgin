library verilog;
use verilog.vl_types.all;
entity simulation_assignment_task_1 is
end simulation_assignment_task_1;
