library verilog;
use verilog.vl_types.all;
entity simualtion_assignment_task_5 is
end simualtion_assignment_task_5;
