library verilog;
use verilog.vl_types.all;
entity simulation_assignment_task_2 is
end simulation_assignment_task_2;
