library verilog;
use verilog.vl_types.all;
entity simulation_task_3 is
end simulation_task_3;
