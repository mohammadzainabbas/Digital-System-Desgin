library verilog;
use verilog.vl_types.all;
entity stimulus_Q4_Assignment2 is
end stimulus_Q4_Assignment2;
