library verilog;
use verilog.vl_types.all;
entity Task_1 is
    port(
        in1             : in     vl_logic;
        in2             : in     vl_logic;
        eq              : out    vl_logic
    );
end Task_1;
