library verilog;
use verilog.vl_types.all;
entity task1 is
    port(
        b1              : in     vl_logic;
        b2              : in     vl_logic;
        b3              : in     vl_logic;
        b4              : in     vl_logic;
        g1              : out    vl_logic;
        g2              : out    vl_logic;
        g3              : out    vl_logic;
        g4              : out    vl_logic
    );
end task1;
