library verilog;
use verilog.vl_types.all;
entity simulation_task_1 is
end simulation_task_1;
