library verilog;
use verilog.vl_types.all;
entity stim is
end stim;
